library verilog;
use verilog.vl_types.all;
entity trcut_tb is
end trcut_tb;
