library verilog;
use verilog.vl_types.all;
entity SDFFtb is
end SDFFtb;
