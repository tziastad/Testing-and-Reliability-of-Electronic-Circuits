library verilog;
use verilog.vl_types.all;
entity TRCUTwithLFSR is
    port(
        CLK             : in     vl_logic;
        SE              : in     vl_logic;
        SO              : out    vl_logic
    );
end TRCUTwithLFSR;
