library verilog;
use verilog.vl_types.all;
entity MyDFFtb is
end MyDFFtb;
