library verilog;
use verilog.vl_types.all;
entity tap_controller_tb is
end tap_controller_tb;
