library verilog;
use verilog.vl_types.all;
entity TRCUTwithMISR_tb is
end TRCUTwithMISR_tb;
