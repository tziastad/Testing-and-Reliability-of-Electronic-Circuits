library verilog;
use verilog.vl_types.all;
entity comb_logic_tb is
end comb_logic_tb;
